module	tb_mux2to1	;

reg	in0	;
reg	in1	;
reg	sel	;
